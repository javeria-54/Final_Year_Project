module controller (
    input  logic clk,
    input  logic reset,
    input  logic start,          
    output logic done           
);

endmodule